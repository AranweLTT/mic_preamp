** Profile: "cascade-total_tdh"  [ G:\workspace\capture\projet_ampli_microphone-pspicefiles\cascade\total_tdh.sim ] 

** Creating circuit file "total_tdh.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of Z:\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 100us 10n 
.FOUR 5k 20 V([VS5]) 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\cascade.net" 


.END
