** Profile: "ampli_diff_5V-diff_simu_gain"  [ D:\lorenzo\projet_ampli_microphone-PSpiceFiles\ampli_diff_5V\diff_simu_gain.sim ] 

** Creating circuit file "diff_simu_gain.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of Z:\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 10Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\ampli_diff_5V.net" 


.END
