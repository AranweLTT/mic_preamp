** Profile: "cascade-total_tdh"  [ D:\lorenzo\capture\projet_ampli_microphone-pspicefiles\cascade\total_tdh.sim ] 

** Creating circuit file "total_tdh.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of Z:\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 100us 5n 
.FOUR 5k 20 V([VS4]) V([VS3]) V([VS2]) V([VS1]) 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\cascade.net" 


.END
